LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY T11_StdLogicVector_Tb IS
END T11_StdLogicVector_Tb;


ARCHITECTURE T11_StdLogicVector_Arch of T11_StdLogicVector_Tb IS
	SIGNAL Slv1: STD_LOGIC_VECTOR(7  DOWNTO 0);
	SIGNAL Slv2: STD_LOGIC_VECTOR(7  DOWNTO 0) := (OTHERS => '0');
	SIGNAL Slv3: STD_LOGIC_VECTOR(7  DOWNTO 0) := (OTHERS => '1');
	SIGNAL Slv4: STD_LOGIC_VECTOR(7  DOWNTO 0) := X"AA";
	SIGNAL Slv5: STD_LOGIC_VECTOR(0  TO 7)     := "10101010";
	SIGNAL Slv6: STD_LOGIC_VECTOR(7  DOWNTO 0) := "00000001";
BEGIN 

	-- Shift Register
	PROCESS IS
	BEGIN 
		
		WAIT FOR 10 NS;
		--FOR i IN 7 DOWNTO 1 loop
		FOR i IN Slv6'LEFT DOWNTO Slv6'RIGHT + 1 loop
			Slv6(i) <= Slv6(i-1);
		END LOOP;
		Slv6(Slv6'RIGHT) <= Slv6(Slv6'LEFT);
 	END PROCESS;



END T11_StdLogicVector_Arch;